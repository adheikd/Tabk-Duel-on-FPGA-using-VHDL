library ieee;
use ieee.std_logic_1164.all;

package tank_const IS
    constant t_size   : INTEGER := 30;
    constant c_length : INTEGER := 0;
    constant c_width  : INTEGER := 14;
    constant b_width  : INTEGER := 5;
    constant bullet_travel : INTEGER := 8;
end package tank_const;
package BODY tank_const is
end package BODY tank_const;